`timescale 1ns / 1ps
module SEG_LUT(
   input[3:0] Q0,
   input[3:0] Q1,
   input[3:0] Q2,
   input[3:0] Q3,
   input[3:0] Q4,  
   input[3:0] Q5,
   input[2:0] sel,
   output reg[5:0] dig,
   output reg[7:0] smg
   );
   always @(*)
   begin 
	case(sel)
		3'd0: 
       begin 
        dig = 6'b011111;
         case(Q0)
		4'd0:smg = 8'b0111_1110;//"0"  8'b1000_0001  8'b0111_1110
		4'd1:smg = 8'b0011_0000;//"1"  8'b1100_1111  8'b0011_0000
		4'd2:smg = 8'b0110_1101;//"2"  8'b1001_0010  8'b0110_1101
		4'd3:smg = 8'b0111_1001;//"3"  8'b1000_0110  8'b0111_1001
		4'd4:smg = 8'b0011_0011;//"4"  8'b1100_1100  8'b0011_0011
		4'd5:smg = 8'b0101_1011;//"5"  8'b1010_0100  8'b0101_1011
		4'd6:smg = 8'b0101_1111;//"6"  8'b1010_0000  8'b0101_1111
		4'd7:smg = 8'b0111_0000;//"7"  8'b1000_1111  8'b0111_0000
		4'd8:smg = 8'b0111_1111;//"8"  8'b1000_0000  8'b0111_1111
		4'd9:smg = 8'b0111_1011;//"9"  8'b1000_0100  8'b0111_1011
		default:smg = 8'b1111_1111;	
	endcase
       end
		3'd1: 
       begin 
        dig = 6'b101111;
        case(Q1)
		4'd0:smg = 8'b0111_1110;//"0"  8'b1000_0001  8'b0111_1110
		4'd1:smg = 8'b0011_0000;//"1"  8'b1100_1111  8'b0011_0000
		4'd2:smg = 8'b0110_1101;//"2"  8'b1001_0010  8'b0110_1101
		4'd3:smg = 8'b0111_1001;//"3"  8'b1000_0110  8'b0111_1001
		4'd4:smg = 8'b0011_0011;//"4"  8'b1100_1100  8'b0011_0011
		4'd5:smg = 8'b0101_1011;//"5"  8'b1010_0100  8'b0101_1011
		4'd6:smg = 8'b0101_1111;//"6"  8'b1010_0000  8'b0101_1111
		4'd7:smg = 8'b0111_0000;//"7"  8'b1000_1111  8'b0111_0000
		4'd8:smg = 8'b0111_1111;//"8"  8'b1000_0000  8'b0111_1111
		4'd9:smg = 8'b0111_1011;//"9"  8'b1000_0100  8'b0111_1011
		default:smg = 8'b1111_1111;		
	endcase
       end 
		3'd2: 
       begin 
        dig = 6'b110111;
        case(Q2)
		4'd0:smg = 8'b1111_1110;//"0"  8'b1000_0001  8'b0111_1110
		4'd1:smg = 8'b1011_0000;//"1"  8'b1100_1111  8'b0011_0000
		4'd2:smg = 8'b1110_1101;//"2"  8'b1001_0010  8'b0110_1101
		4'd3:smg = 8'b1111_1001;//"3"  8'b1000_0110  8'b0111_1001
		4'd4:smg = 8'b1011_0011;//"4"  8'b1100_1100  8'b0011_0011
		4'd5:smg = 8'b1101_1011;//"5"  8'b1010_0100  8'b0101_1011
		4'd6:smg = 8'b1101_1111;//"6"  8'b1010_0000  8'b0101_1111
		4'd7:smg = 8'b1111_0000;//"7"  8'b1000_1111  8'b0111_0000
		4'd8:smg = 8'b1111_1111;//"8"  8'b1000_0000  8'b0111_1111
		4'd9:smg = 8'b1111_1011;//"9"  8'b1000_0100  8'b0111_1011
		default:smg = 8'b1111_1111;		
	endcase
       end 
		3'd3: 
       begin 
        dig = 6'b111011;
        case(Q3)
		4'd0:smg = 8'b0111_1110;//"0"  8'b1000_0001  8'b0111_1110
		4'd1:smg = 8'b0011_0000;//"1"  8'b1100_1111  8'b0011_0000
		4'd2:smg = 8'b0110_1101;//"2"  8'b1001_0010  8'b0110_1101
		4'd3:smg = 8'b0111_1001;//"3"  8'b1000_0110  8'b0111_1001
		4'd4:smg = 8'b0011_0011;//"4"  8'b1100_1100  8'b0011_0011
		4'd5:smg = 8'b0101_1011;//"5"  8'b1010_0100  8'b0101_1011
		4'd6:smg = 8'b0101_1111;//"6"  8'b1010_0000  8'b0101_1111
		4'd7:smg = 8'b0111_0000;//"7"  8'b1000_1111  8'b0111_0000
		4'd8:smg = 8'b0111_1111;//"8"  8'b1000_0000  8'b0111_1111
		4'd9:smg = 8'b0111_1011;//"9"  8'b1000_0100  8'b0111_1011
		default:smg = 8'b1111_1111;	
	endcase
      end
		3'd4: 
       begin 
        dig = 6'b111101;
         case(Q4)
		4'd0:smg = 8'b1111_1110;//"0"  8'b1000_0001  8'b0111_1110
		4'd1:smg = 8'b1011_0000;//"1"  8'b1100_1111  8'b0011_0000
		4'd2:smg = 8'b1110_1101;//"2"  8'b1001_0010  8'b0110_1101
		4'd3:smg = 8'b1111_1001;//"3"  8'b1000_0110  8'b0111_1001
		4'd4:smg = 8'b1011_0011;//"4"  8'b1100_1100  8'b0011_0011
		4'd5:smg = 8'b1101_1011;//"5"  8'b1010_0100  8'b0101_1011
		4'd6:smg = 8'b1101_1111;//"6"  8'b1010_0000  8'b0101_1111
		4'd7:smg = 8'b1111_0000;//"7"  8'b1000_1111  8'b0111_0000
		4'd8:smg = 8'b1111_1111;//"8"  8'b1000_0000  8'b0111_1111
		4'd9:smg = 8'b1111_1011;//"9"  8'b1000_0100  8'b0111_1011
		default:smg = 8'b1111_1111;		
	endcase
       end
		3'd5: 
       begin 
        dig = 6'b111110;
        case(Q5)
		4'd0:smg = 8'b0111_1110;//"0"  8'b1000_0001  8'b0111_1110
		4'd1:smg = 8'b0011_0000;//"1"  8'b1100_1111  8'b0011_0000
		4'd2:smg = 8'b0110_1101;//"2"  8'b1001_0010  8'b0110_1101
		4'd3:smg = 8'b0111_1001;//"3"  8'b1000_0110  8'b0111_1001
		4'd4:smg = 8'b0011_0011;//"4"  8'b1100_1100  8'b0011_0011
		4'd5:smg = 8'b0101_1011;//"5"  8'b1010_0100  8'b0101_1011
		4'd6:smg = 8'b0101_1111;//"6"  8'b1010_0000  8'b0101_1111
		4'd7:smg = 8'b0111_0000;//"7"  8'b1000_1111  8'b0111_0000
		4'd8:smg = 8'b0111_1111;//"8"  8'b1000_0000  8'b0111_1111
		4'd9:smg = 8'b0111_1011;//"9"  8'b1000_0100  8'b0111_1011
		default:smg = 8'b1111_1111;		
	endcase
       end 
       default: dig = 6'b111111;
	endcase
   end
endmodule
